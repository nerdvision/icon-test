vhdl test file
